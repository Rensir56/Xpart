`timescale 1ns/1ps
module MaskGen(
    input  [2:0] memdata_width,
    input [2:0] alu_out,
    input [63:0] rs2_data,
    output reg [7:0] mask_out,
    output reg [63:0] rw_wdata
);

    always@(*) begin
        case(memdata_width)
            3'b000:begin
                mask_out=8'b00000000;
                rw_wdata=rs2_data;
            end
            3'b001:begin
                mask_out=8'b11111111;
                rw_wdata=rs2_data;
            end
            3'b010:begin
                case(alu_out[2])
                    1'b0:begin 
                        mask_out=8'b00001111;
                        rw_wdata=rs2_data;
                    end
                    1'b1:begin
                        mask_out=8'b11110000;
                        rw_wdata=rs2_data<<32;
                    end
                endcase
            end
            3'b011:begin
                case(alu_out[2:1])
                    2'b00:begin
                        mask_out=8'b00000011;
                        rw_wdata=rs2_data;
                    end
                    2'b01:begin
                        mask_out=8'b00001100;
                        rw_wdata=rs2_data<<16;
                    end
                    2'b10:begin
                        mask_out=8'b00110000;
                        rw_wdata=rs2_data<<32;
                    end
                    2'b11:begin
                        mask_out=8'b11000000;
                        rw_wdata=rs2_data<<48;
                    end
                endcase
            end
            3'b100:begin
                case(alu_out[2:0])
                    3'b000:begin
                        mask_out=8'b00000001;
                        rw_wdata=rs2_data;
                    end
                    3'b001:begin
                        mask_out=8'b00000010;
                        rw_wdata=rs2_data<<8;
                    end
                    3'b010:begin
                        mask_out=8'b00000100;
                        rw_wdata=rs2_data<<16;
                    end
                    3'b011:begin
                        mask_out=8'b00001000;
                        rw_wdata=rs2_data<<24;
                    end
                    3'b100:begin
                        mask_out=8'b00010000;
                        rw_wdata=rs2_data<<32;
                    end
                    3'b101:begin
                        mask_out=8'b00100000;
                        rw_wdata=rs2_data<<40;
                    end
                    3'b110:begin
                        mask_out=8'b01000000;
                        rw_wdata=rs2_data<<48;
                    end
                    3'b111:begin
                        mask_out=8'b10000000;
                        rw_wdata=rs2_data<<56;
                    end
                endcase
            end
            3'b101:begin
                case(alu_out[2])
                    1'b0:begin 
                        mask_out=8'b00001111;
                        rw_wdata=rs2_data;
                    end
                    1'b1:begin
                        mask_out=8'b11110000;
                        rw_wdata=rs2_data<<32;
                    end
                endcase
            end
            3'b110:begin
                case(alu_out[2:1])
                    2'b00:begin
                        mask_out=8'b00000011;
                        rw_wdata=rs2_data;
                    end
                    2'b01:begin
                        mask_out=8'b00001100;
                        rw_wdata=rs2_data<<16;
                    end
                    2'b10:begin
                        mask_out=8'b00110000;
                        rw_wdata=rs2_data<<32;
                    end
                    2'b11:begin
                        mask_out=8'b11000000;
                        rw_wdata=rs2_data<<48;
                    end
                endcase
            end
            3'b111:begin
                case(alu_out)
                    3'b000:begin
                        mask_out=8'b00000001;
                        rw_wdata=rs2_data;
                    end
                    3'b001:begin
                        mask_out=8'b00000010;
                        rw_wdata=rs2_data<<8;
                    end
                    3'b010:begin
                        mask_out=8'b00000100;
                        rw_wdata=rs2_data<<16;
                    end
                    3'b011:begin
                        mask_out=8'b00001000;
                        rw_wdata=rs2_data<<24;
                    end
                    3'b100:begin
                        mask_out=8'b00010000;
                        rw_wdata=rs2_data<<32;
                    end
                    3'b101:begin
                        mask_out=8'b00100000;
                        rw_wdata=rs2_data<<40;
                    end
                    3'b110:begin
                        mask_out=8'b01000000;
                        rw_wdata=rs2_data<<48;
                    end
                    3'b111:begin
                        mask_out=8'b10000000;
                        rw_wdata=rs2_data<<56;
                    end
                endcase
            end
        endcase
    end
endmodule